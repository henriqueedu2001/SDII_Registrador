module processor(

);
    
endmodule