module register_file(
    input [7:0] data_input,
    output [7:0] data_output
);
    /* (TODO) */
    assign data_output = data_input;
endmodule