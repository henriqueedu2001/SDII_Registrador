`timescale 1ns/1ps

/* módulo de teste para a rom */
module test_processor #(parameter WORDSIZE = 64, parameter SIZE = 32);
    
endmodule
