module data_memory(
    input [7:0] data_input,
    output [7:0] data_output
);
    assign data_output = data_input;
endmodule